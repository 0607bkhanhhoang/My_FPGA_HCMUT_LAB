library verilog;
use verilog.vl_types.all;
entity sine_wave_generator_vlg_vec_tst is
end sine_wave_generator_vlg_vec_tst;
